library verilog;
use verilog.vl_types.all;
entity MEM_4x3_vlg_vec_tst is
end MEM_4x3_vlg_vec_tst;
