library verilog;
use verilog.vl_types.all;
entity Memoria4x3_vlg_vec_tst is
end Memoria4x3_vlg_vec_tst;
